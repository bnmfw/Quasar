* Analise MC
.param phig_var_p = 4.712547428000001
.param phig_var_n = 4.357688986666666