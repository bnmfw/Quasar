* *       NGLibraryCreator, v2009.07-HR28-2009-07-08 - build 0907160200        *
* *                                                                            *
* ******************************************************************************
* 
* 
*

.GLOBAL VDD
.GLOBAL VSS

********************************************************************************
*                                                                              *
* Cellname:   DFF_X2.                                                          
* Technology: 7nm ASAP
* Format:     Default.                                                         
********************************************************************************
*******.include 7nm_FF.pm

.SUBCKT DFF CK D Q QN VDD VSS //era DFF_X1, eu tirei pq n pode ter X no meu roteiro :)
M_MN2 ci cni VSS VSS nmos_rvt nfin = 1
M_MN6 VSS z4 z6 VSS nmos_rvt nfin = 1
M_MN7 z3 ci z6 VSS nmos_rvt nfin = 1
M_MN4 z2 cni z3 VSS nmos_rvt nfin = 1
M_MN3 z2 D VSS VSS nmos_rvt nfin = 1
M_MN5 z4 z3 VSS VSS nmos_rvt nfin = 1
M_MN1 VSS CK cni VSS nmos_rvt nfin = 1
M_MN8 z12 z3 VSS VSS nmos_rvt nfin = 1
M_MN9 z9 ci z12 VSS nmos_rvt nfin = 1
M_MN12 z9 cni z8 VSS nmos_rvt nfin = 1
M_MN11 z8 z10 VSS VSS nmos_rvt nfin = 1
M_MN10 VSS z9 z10 VSS nmos_rvt nfin = 1
M_MN13 VSS z10 Q VSS nmos_rvt nfin = 1
M_MN14 QN z9 VSS VSS nmos_rvt nfin = 1
M_MP2 ci cni VDD VDD pmos_rvt nfin = 1
M_MP6 VDD z4 z1 VDD pmos_rvt nfin = 1
M_MP7 z1 cni z3 VDD pmos_rvt nfin = 1
M_MP4 z3 ci z5 VDD pmos_rvt nfin = 1
M_MP3 z5 D VDD VDD pmos_rvt nfin = 1
M_MP5 z4 z3 VDD VDD pmos_rvt nfin = 1
M_MP1 VDD CK cni VDD pmos_rvt nfin = 1
M_MP8 z7 z3 VDD VDD pmos_rvt nfin = 1
M_MP9 z9 cni z7 VDD pmos_rvt nfin = 1
M_MP12 z9 ci z11 VDD pmos_rvt nfin = 1
M_MP11 z11 z10 VDD VDD pmos_rvt nfin = 1
M_MP10 VDD z9 z10 VDD pmos_rvt nfin = 1
M_MP13 VDD z10 Q VDD pmos_rvt nfin = 1
M_MP14 QN z9 VDD VDD pmos_rvt nfin = 1
.ENDS 

********************************************************************************
*
* END
*
********************************************************************************

