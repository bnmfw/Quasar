Nand Parsing Test

****** Dispositivos Lógicos ******

.include ../include.cir

****** HGSPICE ******

.option measform = 3
.option post = 2

****** Circuito ******

Xinva1 vcc vss a fa NOT
Xinva2 vcc vss fa ta NOT
Xinvb1 vcc vss b fb NOT
Xinvb2 vcc vss fb tb NOT

****** START QUASAR ******

Mp11 vdd ta g1 ta PMOS_RVT nfin=3
Mp12 vdd tb g1 tb PMOS_RVT nfin=3
Mn11 g1 ta i1 ta NMOS_RVT nfin=3
Mn12 i1 tb vss tb NMOS_RVT nfin=3

****** END QUASAR ******

//Representação de um circuito pós benchmark
xff1 clk g1 q1 nq1 vcc vss DFF
xinv11 vcc vss q1 nnq1 NOT

************
.end