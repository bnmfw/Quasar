Benchmark C17 V0

****** Dispositivos Lógicos ******

.include dis/logica.cir
.include dis/DFF.cir
.include mc.cir

****** HGSPICE ******

.option measform = 3
.option post = 0

****** Fontes de Tensão Geral ******

.include vdd.cir

****** Fontes de Sinal ******

.include fontes.cir

****** SETs ******

.include SETs.cir

****** Circuito ******

Xinva1 vcc gnd a fa NOT
Xinva2 vcc gnd fa ta NOT
Xinvb1 vcc gnd b fb NOT
Xinvb2 vcc gnd fb tb NOT

Mp11 vdd ta g1 ta PMOS_RVT nfin=3
Mp12 vdd tb g1 tb PMOS_RVT nfin=3
Mn11 g1 ta i1 ta NMOS_RVT nfin=3
Mn12 i1 tb gnd tb NMOS_RVT nfin=3

Vmeasg1 g1 m1 0

//Representação de um circuito pós benchmark
xff1 clk m1 q1 nq1 vcc gnd DFF
xinv11 vcc gnd q1 nnq1 NOT

****** Controle ******

.include largura_pulso.cir
.include atraso.cir
.include monte_carlo.cir

************
.end
