Nor

****** Dispositivos Lógicos ******

.include ../../include.cir

****** Circuito ******

Mp1 vdd a i1 vdd PMOS W=140n L=32n
Mp2 i1 b g1 vdd PMOS W=140n L=32n
Mn1 g1 a gnd gnd NMOS W=70n L=32n
Mn2 g1 b gnd gnd NMOS W=70n L=32n

Mp3 vdd g1 ng1 vdd PMOS W=140n L=32n    
Mn3 ng1 g1 gnd gnd NMOS W=70n L=32n

****** END QUASAR ******

************
.end