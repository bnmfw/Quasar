Nand

****** Dispositivos Lógicos ******

.include ../include.cir

****** HGSPICE ******

.option measform = 3
.option post = 0

****** Circuito ******

Mp1 vdd a fa vdd PMOS_RVT nfin=3
Mn1 fa a gnd gnd NMOS_RVT nfin=3
Mp2 vdd b fb vdd PMOS_RVT nfin=3
Mn2 fb b gnd gnd NMOS_RVT nfin=3

Mp3 vdd fa ta vdd PMOS_RVT nfin=3
Mn3 ta fa gnd gnd NMOS_RVT nfin=3
Mp4 vdd fb tb vdd PMOS_RVT nfin=3
Mn4 tb fb gnd gnd NMOS_RVT nfin=3

Mp11 vdd ta g1 vdd PMOS_RVT nfin=3
Mp12 vdd tb g1 vdd PMOS_RVT nfin=3
Mn11 g1 ta i1 gnd NMOS_RVT nfin=3
Mn12 i1 tb gnd gnd NMOS_RVT nfin=3

//Representação de um circuito pós benchmark
xff1 clk g1 q1 nq1 vcc gnd DFF
xinv11 vcc gnd q1 nnq1 NOT

************
.end