.include ../../include.cir
.option measform = 3
.option post = 0

* DECLARANDO O CIRCUITO
Mp0	vdd	SELECT	n1	vdd	PMOS w=105n l=32n
Mn0 	n1 	SELECT 	gnd 	gnd	NMOS w=70n  l=32n

Mp1 	vdd 	n1 	x1 	vdd	PMOS w=105n l=32n
Mp2 	vdd 	A 	x1 	vdd 	PMOS w=105n l=32n
Mn1 	x1 	n1 	n2 	gnd	NMOS w=140n l=32n
Mn2	n2	A	gnd	gnd	NMOS w=140n l=32n

Mp3 	vdd 	SELECT 	x2 	vdd	PMOS w=105n l=32n
Mp4 	vdd 	B 	x2 	vdd 	PMOS w=105n l=32n
Mn3 	x2 	SELECT 	n3 	gnd	NMOS w=140n l=32n
Mn4	n3	B	gnd	gnd	NMOS w=140n l=32n

Mp5 	vdd 	x2 	out 	vdd	PMOS w=105n l=32n
Mp6 	vdd 	x1 	out 	vdd 	PMOS w=105n l=32n
Mn5 	out 	x1 	n4 	gnd	NMOS w=140n l=32n
Mn6	n4	x2	gnd	gnd	NMOS w=140n l=32n

MpC1E1	vdd	inA	a2	vdd	PMOS  w=105n  l=32n
MnC1E1	a2	inA	gnd	gnd	NMOS  w=70n   l=32n

MpC2E1	vdd	a2	A	vdd	PMOS  w=105n  l=32n
MnC2E1	A	a2	gnd	gnd	NMOS  w=70n   l=32n

MpC1E2	vdd	inB	b2	vdd	PMOS  w=105n  l=32n
MnC1E2	b2	inB	gnd	gnd	NMOS  w=70n   l=32n

MpC2E2	vdd	b2	B	vdd	PMOS  w=105n  l=32n
MnC2E2	B	b2	gnd	gnd	NMOS  w=70n   l=32n

MpC1E3	vdd	inSel	sel2	vdd	PMOS  w=105n  l=32n
MnC1E3	sel2	inSel	gnd	gnd	NMOS  w=70n   l=32n

MpC2E3	vdd	sel2	SELECT	vdd	PMOS  w=105n  l=32n
MnC2E3	SELECT	sel2	gnd	gnd	NMOS  w=70n   l=32n

Cload	out	gnd	100f

.end