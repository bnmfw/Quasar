**** Unidades de memória ****

**** Dispositivos logicos ****

.include logica.cir
.include multiplex.cir

**** Subcircuito FLIP FLOP JK ****

.subckt FFJK vp vm j k clk q nq
c1 clk clkt 0.1n
r1 clkt gnd 0.5
xnand1 vp vm j clkt 1 NAND
xnand2 vp vm k clkt 2 NAND
xnand3 vp vm 1 nq q NAND
xnand4 vp vm 2 q nq NAND
.ends

**** Subcircuito FLIP FLOP T ****

.subckt FFT vp vm t clk q nq
c1 clk clkt 0.1n
r1 clkt gnd 0.5
xnand1 vp vm t clkt nq 1 NAND3
xnand2 vp vm t clkt q 2 NAND3
xnand3 vp vm 1 nq q NAND
xnand4 vp vm 2 q nq NAND
*Cload1  q gnd 0.5
*Cload2 nq vdd 0.5
.ends

**** Subcircuito FLIP FLOP D ****

* 11 pares CMOS *
.subckt FFD vp vm d clk q nq
xnot1 vp vm clk nclk NOT
xlatch1 vp vm d nclk qm 1 LTD
xlatch2 vp vm qm clk q 2 LTD
.ends

**** Subcircuito LATCH JK ****

.subckt LATCHJK vp vm j k clk q nq
xnand1 vp vm j clk 1 NAND
xnand2 vp vm k clk 2 NAND
xnand3 vp vm 1 nq q NAND
xnand4 vp vm 2 q nq NAND
.ends 

**** Subcircuito LATCH D ****

* 5 pares CMOS *
.subckt LTD vp vm d clk q nq
xmux vp vm d 1 clk q MUX1
xnot1 vp vm q nq NOT
xnot2 vp vm nq 1 NOT
.ends

**** Subcircuito LATCH T ****

.subckt LATCHT vp vm t clk q nq
xnand1 vp vm t clk q 1 NAND3
xnand2 vp vm t clk nq 2 NAND3
xnand3 vp vm 1 nq q NAND
xnand4 vp vm 2 q nq NAND
.ends 

.end

