* Analise MC
.param phig_var_p = 4.596727418
.param phig_var_n = 4.3187854733333335