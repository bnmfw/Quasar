Arquivo para testar minhas bibliotecas
** DAAABBBBB*** 


****** Finfets ******

.include logica.cir

****** Fontes de Tensão Geral ******

Vvdd vdd gnd 0.7 

****** Fontes de Sinal ******

Va a gnd PULSE(0 0.9  5n 0.01n 0.01n  5n  10n)
Vb b gnd PULSE(0 0.9 10n 0.01n 0.01n 10n  20n)
Vc c gnd PULSE(0 0.9 20n 0.01n 0.01n 20n  40n)
Vd d gnd PULSE(0 0.9 40n 0.01n 0.01n 40n  80n)
Ve e gnd PULSE(0 0.9 80n 0.01n 0.01n 80n 160n)

****** Circuito ******

xnot vdd gnd a s NOT
ca s gnd 1f

****** Controle ******

.tran 10ps 160ns
.plot v(a) v(s)
.option measform = 3 //gera a saída em .csv
.option post = 2 //permite o uso do cscope

*.meas tran FallA TRIG v(a) val='0.35' rise=1 TARG v(s) val='0.35' fall=1
*.meas tran RiseA TRIG v(a) val='0.35' fall=1 TARG v(s) val='0.35' rise=1
*.meas tran Corr INTEG i(Vvdd) from=0 to=25n

****************
.end
