Nor Parsing Test

****** Dispositivos Lógicos ******

.include ../../include.cir

****** Circuito ******

Xinva1 vcc gnd a fa NOT
Xinva2 vcc gnd fa ta NOT
Xinvb1 vcc gnd b fb NOT
Xinvb2 vcc gnd fb tb NOT

****** START QUASAR ******

Mp51 vdd ta i1 ta PMOS_RVT nfin=3
Mp52 i1 tb g1 tb PMOS_RVT nfin=3
Mn51 g1 ta gnd ta NMOS_RVT nfin=3
Mn52 g1 tb gnd tb NMOS_RVT nfin=3

****** END QUASAR ******

//Representação de um circuito pós benchmark
xff1 clk g1 q1 nq1 vcc gnd DFF
xinv11 vcc gnd q1 nnq1 NOT

************
.end