SET Simulation TG

**** Dispositivos Lógicos *******

.include ../include.cir

****** HSPICE ******

.option measform = 3
.option post = 0

**********Circuito******

* ENTRADA inA
MpC1E1	vdd	inA	a2	vdd	PMOS_BULK  w=140n  L=32n
MnC1E1	a2	inA	gnd	gnd	NMOS_BULK  w=70n   L=32n

MpC2E1	vdd	a2	a	vdd	PMOS_BULK  w=140n  L=32n
MnC2E1	a	a2	gnd	gnd	NMOS_BULK  w=70n   L=32n

* ENTRADA inB
MpC1E2	vdd	inB	b2	vdd	PMOS_BULK  w=140n  L=32n
MnC1E2	b2	inB	gnd	gnd	NMOS_BULK  w=70n   L=32n

MpC2E2	vdd	b2	b	vdd	PMOS_BULK  w=140n  L=32n
MnC2E2	b	b2	gnd	gnd	NMOS_BULK  w=70n   L=32n

* ENTRADA inSel
MpC1E3	vdd	inSel	sel2	vdd	PMOS_BULK  w=140n  L=32n
MnC1E3	sel2	inSel	gnd	gnd	NMOS_BULK  w=70n   L=32n

MpC2E3	vdd	sel2	select	vdd	PMOS_BULK  w=140n  L=32n
MnC2E3	select	sel2	gnd	gnd	NMOS_BULK  w=70n   L=32n

Mp0	vdd	select n1 vdd PMOS_BULK w=140n l=32n
Mn0 n1 select gnd gnd NMOS_BULK w=70n l=32n

Mp1 a select out vdd PMOS_BULK w=140n l=32n
Mn1 a n1 out gnd NMOS_BULK w=70n l=32n

Mp2 b n1 out vdd PMOS_BULK w=140n l=32n
Mn2	b select out gnd NMOS_BULK w=70n l=32n


* Fan outs
Mpcs1 vdd out sc1 vdd PMOS_BULK  w=560n  L=32n
Mncs1 sc1 out gnd gnd NMOS_BULK  w=280n  L=32n
Mpcs2 vdd sc1 sc2 vdd PMOS_BULK  w=560n  L=32n
Mncs2 sc2 sc1 gnd gnd NMOS_BULK  w=280n  L=32n

**********************

.end