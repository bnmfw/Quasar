*Arquivo Analise Monte Carlo
.tran 0.01n 4n