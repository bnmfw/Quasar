Xor v5

****** Dispositivos Lógicos ******

.include ../include.cir

****** HGSPICE ******

.option measform = 3
.option post = 0

****** Circuito ******

* Not
Mp1 vdd a na vdd PMOS_RVT nfin=3
Mn1 na a gnd gnd NMOS_RVT nfin=3

* Not
Mp2 vdd b nb vdd PMOS_RVT nfin=3
Mn2 nb b gnd gnd NMOS_RVT nfin=3

Mp3 a b axorb vdd PMOS_RVT nfin=3
Mn3 a nb axorb gnd NMOS_RVT nfin=3

Mp4 na nb axorb vdd PMOS_RVT nfin=3
Mn4 na b axorb gnd NMOS_RVT nfin=3
************
.end