Nand Parsing Test

****** Dispositivos Lógicos ******

.include ../../include.cir

****** START QUASAR ******

Mp11 vdd a g1 vdd PMOS_RVT nfin=3
Mp12 vdd b g1 vdd PMOS_RVT nfin=3
Mn11 g1 a i1 gnd NMOS_RVT nfin=3
Mn12 i1 b gnd gnd NMOS_RVT nfin=3

****** END QUASAR ******

************
.end