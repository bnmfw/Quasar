* Analise MC
.param phig_var_p = gauss(4.8108, 0.05, 3)
.param phig_var_n = gauss(4.372, 0.05, 3)