Xor v1

****** Dispositivos Lógicos ******

.include ../../include.cir

****** Circuito ******

Mp1 vdd a na vdd PMOS_RVT nfin=3
Mn1 na a gnd gnd NMOS_RVT nfin=3

Mp2 vdd b nb vdd PMOS_RVT nfin=3
Mn2 nb b gnd gnd NMOS_RVT nfin=3

Mp3 vdd na i1 vdd PMOS_RVT nfin=3
Mp4 i1 b axorb vdd PMOS_RVT nfin=3
Mp5 vdd a i2 vdd PMOS_RVT nfin=3
Mp6 i2 nb axorb vdd PMOS_RVT nfin=3

Mn3 axorb nb i3 gnd NMOS_RVT nfin=3
Mn4 i3 na gnd gnd NMOS_RVT nfin=3
Mn5 axorb b i4 gnd NMOS_RVT nfin=3
Mn6 i4 a gnd gnd NMOS_RVT nfin=3
************
.end