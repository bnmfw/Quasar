Nand

****** Dispositivos Lógicos ******

.include ../../include.cir

****** HGSPICE ******

.option measform = 3
.option post = 0

****** Circuito ******

Mp11 vdd a g1 vdd PMOS w=140n L=32n
Mp12 vdd b g1 vdd PMOS w=140n L=32n
Mn11 g1 a i1 gnd NMOS w=70n L=32n
Mn12 i1 b gnd gnd NMOS w=70n L=32n

************
.end