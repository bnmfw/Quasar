Nand Parsing Test

****** Dispositivos Lógicos ******

.include ../include.cir

****** HGSPICE ******

.option measform = 3
.option post = 2

****** START QUASAR ******

Mp11 vdd a g1 vdd PMOS_RVT nfin=3
Mp12 vdd b g1 vdd PMOS_RVT nfin=3
Mn11 g1 a i1 vss NMOS_RVT nfin=3
Mn12 i1 b vss vss NMOS_RVT nfin=3

****** END QUASAR ******

//Representação de um circuito pós benchmark
xff1 clk g1 q1 nq1 vcc vss DFF
xinv11 vcc vss q1 nnq1 NOT

************
.end