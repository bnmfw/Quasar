Nor3

****** Dispositivos Lógicos ******

.include ../../include.cir

****** HGSPICE ******

.option measform = 3
.option post = 0

****** Circuito ******

Mp1 vdd a i1 vdd PMOS_RVT nfin=3
Mp2 i1 b i2 vdd PMOS_RVT nfin=3
Mp3 i2 c g1 vdd PMOS_RVT nfin=3
Mn1 g1 a gnd gnd NMOS_RVT nfin=3
Mn2 g1 b gnd gnd NMOS_RVT nfin=3
Mn3 g1 c gnd gnd NMOS_RVT nfin=3

Mp4 vdd g1 ng1 vdd PMOS_RVT nfin=4
Mn4 ng1 g1 gnd gnd NMOS_RVT nfin=4

************
.end