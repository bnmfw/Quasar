**** Operadores matemáticos usando cmos ****

**** Finfets ****

.include 7nm_FF.pm

**** Dispositivos logicos ****

.include logica.cir

**** Subcircuito Half adder ****

.subckt HADD vp vm a b sum cout
xand1 vp vm a b cout AND
xxor vp vm a b sum XOR
*CloadS sum gnd 10f
*CloadC cout gnd 10f
.ends

**** Subcircuito Full adder ****

.subckt FADD vp vm a b cin sum cout
Mp1 vp a 1 a PMOS_RVT nfin=3
Mp2 1 b ncout b PMOS_RVT nfin=3

Mn1 ncout a 2 a NMOS_RVT nfin=3
Mn2 2 b vm b NMOS_RVT nfin=3

Mp3 vp a 3 a PMOS_RVT nfin=3
Mp4 vp b 3 b PMOS_RVT nfin=3
Mp5 3 cin ncout cin PMOS_RVT nfin=3

Mn3 ncout cin 4 cin NMOS_RVT nfin=3
Mn4 4 a vm a NMOS_RVT nfin=3
Mn5 4 b vm b NMOS_RVT nfin=3

Mp6 vp a 5 a PMOS_RVT nfin=3
Mp7 vp b 5 b PMOS_RVT nfin=3
Mp8 vp cin 5 cin PMOS_RVT nfin=3
Mp9 5 ncout nsum ncout PMOS_RVT nfin=3

Mn6 nsum ncout 6 ncout NMOS_RVT nfin=3
Mn7 6 a vm a NMOS_RVT nfin=3n
Mn8 6 b vm a NMOS_RVT nfin=3
Mn9 6 cin vm cin NMOS_RVT nfin=3

Mp10 vp a 7 a PMOS_RVT nfin=3
Mp11 7 b 8 b PMOS_RVT nfin=3
Mp12 8 cin nsum cin PMOS_RVT nfin=3

Mn10 nsum a 9 a NMOS_RVT nfin=3
Mn11 9 b 10 b NMOS_RVT nfin=3
Mn12 10 cin vm cin NMOS_RVT nfin=3

Mp13 vp nsum sum nsum PMOS_RVT nfin=3
Mn13 sum nsum vm nsum NMOS_RVT nfin=3
Mp14 vp ncout cout ncout PMOS_RVT nfin=3
Mn14 cout ncout vm ncout NMOS_RVT nfin=3

.ends

**** Subcircuito Somador 4 bits ****

.subckt SOM4 vp vm a0 a1 a2 a3 b0 b1 b2 b3 s0 s1 s2 s3 cout
xhadd vp vm a0 b0 s0 c0 HADD
xfadd1 vp vm a1 b1 c0 s1 c1 FADD
xfadd2 vp vm a2 b2 c1 s2 c2 FADD
xfadd3 vp vm a3 b3 c2 s3 cout FADD
.ends
