Xor v5

****** Dispositivos Lógicos ******

.include ../../include.cir

****** HGSPICE ******

.option measform = 3
.option post = 0

****** Circuito ******

Mp11 vdd ta fa vdd PMOS_RVT nfin=3
Mn11 fa ta gnd gnd NMOS_RVT nfin=3
Mp12 vdd fa a vdd PMOS_RVT nfin=3
Mn12 a fa gnd gnd NMOS_RVT nfin=3

Mp13 vdd tb fb vdd PMOS_RVT nfin=3
Mn13 fb tb gnd gnd NMOS_RVT nfin=3
Mp14 vdd fb b vdd PMOS_RVT nfin=3
Mn14 b fb gnd gnd NMOS_RVT nfin=3

* Not
Mp1 vdd a na vdd PMOS_RVT nfin=3
Mn1 na a gnd gnd NMOS_RVT nfin=3

* Not
Mp2 vdd b nb vdd PMOS_RVT nfin=3
Mn2 nb b gnd gnd NMOS_RVT nfin=3

Mp3 a b axorb vdd PMOS_RVT nfin=3
Mn3 a nb axorb gnd NMOS_RVT nfin=3

Mp4 na nb axorb vdd PMOS_RVT nfin=3
Mn4 na b axorb gnd NMOS_RVT nfin=3

Mp15 vdd axorb g1 vdd PMOS_RVT nfin=3
Mn15 g1 axorb gnd gnd NMOS_RVT nfin=3
************
.end