Benchmark C17 V0

****** Dispositivos Lógicos ******

.include ../include.cir

****** HGSPICE ******

.option measform = 3
.option post = 0

****** START QUASAR ******

Mp11 vdd a e1 a PMOS_RVT nfin=3
Mp12 vdd b e1 b PMOS_RVT nfin=3
Mn11 e1 a i1 a NMOS_RVT nfin=3
Mn12 i1 b gnd b NMOS_RVT nfin=3

Mp21 vdd d e2 d PMOS_RVT nfin=3
Mp22 vdd b e2 b PMOS_RVT nfin=3
Mn21 e2 d i2 d NMOS_RVT nfin=3
Mn22 i2 b gnd b NMOS_RVT nfin=3

Mp31 vdd e2 e3 e2 PMOS_RVT nfin=3
Mp32 vdd c e3 c PMOS_RVT nfin=3
Mn31 e3 e2 i3 e2 NMOS_RVT nfin=3
Mn32 i3 c gnd c NMOS_RVT nfin=3

Mp41 vdd e1 g1 e1 PMOS_RVT nfin=3
Mp42 vdd e3 g1 e3 PMOS_RVT nfin=3
Mn41 g1 e1 i4 e1 NMOS_RVT nfin=3
Mn42 i4 e3 gnd e3 NMOS_RVT nfin=3

Mp51 vdd e i5 e PMOS_RVT nfin=3
Mp52 i5 c e4 c PMOS_RVT nfin=3
Mn51 e4 e gnd e NMOS_RVT nfin=3
Mn52 e4 c gnd c NMOS_RVT nfin=3

Mp61 vdd d i62 d PMOS_RVT nfin=3
Mp62 vdd b i62 b PMOS_RVT nfin=3
Mn61 i62 d i61 d NMOS_RVT nfin=3
Mn62 i61 b gnd b NMOS_RVT nfin=3

Mp63 vdd i62 e5 i62 PMOS_RVT nfin=3
Mn63 e5 i62 gnd i62 NMOS_RVT nfin=3

Mp71 vdd e4 i7 e4 PMOS_RVT nfin=3
Mp72 i7 e5 g2 e5 PMOS_RVT nfin=3
Mn71 g2 e4 gnd e4 NMOS_RVT nfin=3
Mn72 g2 e5 gnd e5 NMOS_RVT nfin=3

****** END QUASAR ******

//Representação de um circuito pós benchmark
xff1 clk g1 q1 nq1 vcc gnd DFF
xff2 clk g2 q2 nq2 vcc gnd DFF
xinv11 vcc gnd q1 nnq1 NOT
xinv12 vcc gnd q2 nnq2 NOT  

************
.end
