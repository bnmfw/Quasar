Benchmark C17 V3 (C17_Nand)

****** Dispositivos Logicos ******

.include ../../include.cir

****** HSPICE ******

.option measform = 3
.option post = 0

****** Circuito ******

Mp11 vdd a e1 a PMOS_RVT nfin=3
Mp12 vdd b e1 b PMOS_RVT nfin=3
Mn11 e1 a i1 a NMOS_RVT nfin=3
Mn12 i1 b gnd b NMOS_RVT nfin=3

Mp21 vdd d e2 d PMOS_RVT nfin=3
Mp22 vdd b e2 b PMOS_RVT nfin=3
Mn21 e2 d i2 d NMOS_RVT nfin=3
Mn22 i2 b gnd b NMOS_RVT nfin=3

Mp31 vdd c e3 c PMOS_RVT nfin=3
Mp32 vdd e2 e3 e2 PMOS_RVT nfin=3
Mn31 e3 c i3 c NMOS_RVT nfin=3
Mn32 i3 e2 gnd e2 NMOS_RVT nfin=3

Mp41 vdd e e4 e PMOS_RVT nfin=3
Mp42 vdd e2 e4 e2 PMOS_RVT nfin=3
Mn41 e4 e i4 e NMOS_RVT nfin=3
Mn42 i4 e2 gnd e2 NMOS_RVT nfin=3

Mp51 vdd e1 g1 e1 PMOS_RVT nfin=3
Mp52 vdd e3 g1 e3 PMOS_RVT nfin=3
Mn51 g1 e1 i5 e1 NMOS_RVT nfin=3
Mn52 i5 e3 gnd e3 NMOS_RVT nfin=3

Mp61 vdd e4 g2 e4 PMOS_RVT nfin=3
Mp62 vdd e3 g2 e3 PMOS_RVT nfin=3
Mn61 g2 e4 i6 e4 NMOS_RVT nfin=3
Mn62 i6 e3 gnd e3 NMOS_RVT nfin=3 

************
.end
