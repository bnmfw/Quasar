*mc sweep file
.tran 0.01n 4n