Nor5

****** Dispositivos Lógicos ******

.include ../include.cir

****** HGSPICE ******

.option measform = 3
.option post = 0

****** Circuito ******

Mp1 vdd a i1 vdd PMOS_RVT nfin=3
Mp2 i1 b i2 vdd PMOS_RVT nfin=3
Mp3 i2 c i3 vdd PMOS_RVT nfin=3
Mp4 i3 d i4 vdd PMOS_RVT nfin=3
Mp5 i4 e i5 vdd PMOS_RVT nfin=3
Mp6 i5 f g1 vdd PMOS_RVT nfin=3

Mn1 g1 a gnd gnd NMOS_RVT nfin=3
Mn2 g1 b gnd gnd NMOS_RVT nfin=3
Mn3 g1 c gnd gnd NMOS_RVT nfin=3
Mn4 g1 d gnd gnd NMOS_RVT nfin=3
Mn5 g1 e gnd gnd NMOS_RVT nfin=3
Mn6 g1 f gnd gnd NMOS_RVT nfin=3

Mp10 vdd g1 ng1 vdd PMOS_RVT nfin=4
Mn10 ng1 g1 gnd gnd NMOS_RVT nfin=4

************
.end