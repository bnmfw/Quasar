* Analise MC
.param phig_var_p = 4.7088190580000004
.param phig_var_n = 4.4198005333333334