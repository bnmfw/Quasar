Xor v8

****** Dispositivos Lógicos ******

.include ../../include.cir

****** HGSPICE ******

.option measform = 3
.option post = 0

****** Circuito ******

Mp11 vdd ta fa vdd PMOS_RVT nfin=3
Mn11 fa ta gnd gnd NMOS_RVT nfin=3
Mp12 vdd fa a vdd PMOS_RVT nfin=3
Mn12 a fa gnd gnd NMOS_RVT nfin=3

Mp13 vdd tb fb vdd PMOS_RVT nfin=3
Mn13 fb tb gnd gnd NMOS_RVT nfin=3
Mp14 vdd fb b vdd PMOS_RVT nfin=3
Mn14 b fb gnd gnd NMOS_RVT nfin=3

Mp1 vdd b nb vdd PMOS_RVT nfin=3
Mn1 nb b gnd gnd NMOS_RVT nfin=3

Mp2 a b axorb vdd PMOS_RVT nfin=3
Mn2 a nb axorb gnd NMOS_RVT nfin=3

Mp3 b a axorb vdd PMOS_RVT nfin=3
Mn3 nb a axorb gnd NMOS_RVT nfin=3

************
.end