NAND3

****** Dispositivos Lógicos ******

.include ../include.cir

****** HGSPICE ******

.option measform = 3
.option post = 0

****** Circuito ******

Mp1 vdd a g1 vdd PMOS_BULK w=140n l=32n
Mp2 vdd b g1 vdd PMOS_BULK w=140n l=32n
Mp3 vdd c g1 vdd PMOS_BULK w=140n l=32n
Mn1 g1 a i1 gnd NMOS_BULK w=70n l=32n
Mn2 i1 b i2 gnd NMOS_BULK w=70n l=32n
Mn3 i2 c gnd gnd NMOS_BULK w=70n l=32n

************
.end