Xor v1

****** Dispositivos Lógicos ******

.include ../../include.cir

****** HGSPICE ******

.option measform = 3
.option post = 0

****** Circuito ******

*** FAN IN ****

Mp11 vdd ta fa vdd PMOS_BULK w=140n  L=32n
Mn11 fa ta gnd gnd NMOS_BULK w=70n  L=32n
Mp12 vdd fa a vdd PMOS_BULK w=140n  L=32n
Mn12 a fa gnd gnd NMOS_BULK w=70n  L=32n

Mp13 vdd tb fb vdd PMOS_BULK w=140n  L=32n
Mn13 fb tb gnd gnd NMOS_BULK w=70n  L=32n
Mp14 vdd fb b vdd PMOS_BULK w=140n  L=32n
Mn14 b fb gnd gnd NMOS_BULK w=70n  L=32n

*** CIRCUITO ***

Mp1 vdd a na vdd PMOS_BULK w=140n  L=32n
Mn1 na a gnd gnd NMOS_BULK w=70n  L=32n

Mp2 vdd b nb vdd PMOS_BULK w=140n  L=32n
Mn2 nb b gnd gnd NMOS_BULK w=70n  L=32n

Mp3 vdd na i1 vdd PMOS_BULK w=280n  L=32n
Mp4 i1 b axorb vdd PMOS_BULK w=280n  L=32n
Mp5 vdd a i2 vdd PMOS_BULK w=280n  L=32n
Mp6 i2 nb axorb vdd PMOS_BULK w=280n  L=32n

Mn3 axorb nb i3 gnd NMOS_BULK w=140n  L=32n
Mn4 i3 na gnd gnd NMOS_BULK w=140n  L=32n
Mn5 axorb b i4 gnd NMOS_BULK w=140n  L=32n
Mn6 i4 a gnd gnd NMOS_BULK w=140n  L=32n

*** FAN OUT ***

Mp21 vdd axorb naxorb vdd PMOS_BULK w=560n  L=32n
Mn21 naxorb axorb gnd gnd NMOS_BULK w=280n  L=32n

************
.end