* MUX V19

****** Dispositivos Lógicos ******

.include ../include.cir

****** HSPICE ******

.option measform = 3
.option post = 0

	Mp0	vdd	SELECT	n1	vdd	PMOS w=105n l=32n
	Mn0 	n1 	SELECT 	gnd 	gnd	NMOS w=70n  l=32n

	Mp1 	vdd 	A 	n2 	vdd	PMOS w=105n l=32n
	Mn1 	n2 	A 	gnd 	gnd	NMOS w=70n l=32n

	Mp2 	vdd 	B 	n3 	vdd 	PMOS w=105n l=32n
	Mn2	n3	B	gnd	gnd	NMOS w=70n l=32n

	Mp3	n4	n5	out	vdd	PMOS w=105n l=32n
	Mp4	n6	n4	n5	vdd	PMOS w=105n l=32n
	Mp5	vdd	n4	n6	vdd	PMOS w=105n l=32n
	Mp6	vdd	n5	out	vdd	PMOS w=105n l=32n

	Mn3	A	SELECT	n4	gnd	NMOS w=140n l=32n
	Mn4	B	n1	n4	gnd	NMOS w=140n l=32n
	Mn5 	n2 	SELECT 	n5 	gnd	NMOS w=140n l=32n
	Mn6	n3	n1	n5	gnd	NMOS w=140n l=32n
	Mn7	n6	n4	gnd	gnd	NMOS w=140n l=32n
	Mn8	out	n5	gnd	gnd	NMOS w=140n l=32n

	MpC1E1	vdd	inA	a2	vdd	PMOS  w=105n  l=32n
	MnC1E1	a2	inA	gnd	gnd	NMOS  w=70n   l=32n

	MpC2E1	vdd	a2	A	vdd	PMOS  w=105n  l=32n
	MnC2E1	A	a2	gnd	gnd	NMOS  w=70n   l=32n

	MpC1E2	vdd	inB	b2	vdd	PMOS  w=105n  l=32n
	MnC1E2	b2	inB	gnd	gnd	NMOS  w=70n   l=32n

	MpC2E2	vdd	b2	B	vdd	PMOS  w=105n  l=32n
	MnC2E2	B	b2	gnd	gnd	NMOS  w=70n   l=32n

	MpC1E3	vdd	inSel	sel2	vdd	PMOS  w=105n  l=32n
	MnC1E3	sel2	inSel	gnd	gnd	NMOS  w=70n   l=32n

	MpC2E3	vdd	sel2	SELECT	vdd	PMOS  w=105n  l=32n
	MnC2E3	SELECT	sel2	gnd	gnd	NMOS  w=280n  l=32n

	Mpcs1	vdd	OUT	sc1	vdd	PMOS  w=420n  l=32n
	Mncs1	sc1	OUT	gnd	gnd	NMOS  w=280n  l=32n

	Mpcs2	vdd	sc1	sc2	vdd	PMOS  w=420n  l=32n
	Mncs2	sc2	sc1	gnd	gnd	NMOS  w=280n  l=32n

	.end
