Template

.include ../../include.cir

.option post=2
.option measform=3

*Inversor de entrada do sinal de entrada a1
Mp1 ina a1 vdd vdd pmos_rvt nfin=3
Mn1 gnd a1 ina gnd nmos_rvt nfin=3

*Inversor para a entrada "as" para ficar mais realistico
Mp2 temp_as as vdd vdd pmos_rvt nfin=3
Mn2 gnd as temp_as gnd nmos_rvt nfin=3

Mp3 as_out temp_as vdd vdd pmos_rvt nfin=3
Mn3 gnd temp_as as_out gnd nmos_rvt nfin=3

*Inversor Rad-Hard
Mp4 vdd ina sout vdd pmos_rvt nfin=3
Mn4 sout ina gnd  gnd nmos_rvt nfin=3

Mp5 vdd as_out x vdd pmos_rvt nfin=3
Mn5 x as_out sout gnd nmos_rvt nfin=3

*Inversor de saida do sinal de saida sout
Mp6 s sout vdd vdd pmos_rvt nfin=3
Mn6 gnd sout s gnd nmos_rvt nfin=3

Cload s gnd 1f

.end