Nor

****** Dispositivos Lógicos ******

.include ../include.cir

****** HGSPICE ******

.option measform = 3
.option post = 0

****** Circuito ******

Mp1 vdd a i1 vdd PMOS_RVT nfin=3
Mp2 i1 b g1 vdd PMOS_RVT nfin=3
Mn1 g1 a gnd gnd NMOS_RVT nfin=3
Mn2 g1 b gnd gnd NMOS_RVT nfin=3

Mp3 vdd g1 ng1 vdd PMOS_RVT nfin=4
Mn3 ng1 g1 gnd gnd NMOS_RVT nfin=4

****** END QUASAR ******

//Representação de um circuito pós benchmark
xff1 clk g1 q1 nq1 vcc gnd DFF
xinv11 vcc gnd q1 nnq1 NOT

************
.end